//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This class records instruction_memory transaction information using
//       a covergroup named instruction_memory_transaction_cg.  An instance of this
//       coverage component is instantiated in the uvmf_parameterized_agent
//       if the has_coverage flag is set.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class instruction_memory_transaction_coverage  extends uvm_subscriber #(.T(instruction_memory_transaction ));

  `uvm_component_utils( instruction_memory_transaction_coverage )

  T coverage_trans;

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end
  
  // ****************************************************************************
  covergroup instruction_memory_transaction_cg;
    // pragma uvmf custom covergroup begin
    // UVMF_CHANGE_ME : Add coverage bins, crosses, exclusions, etc. according to coverage needs.
    option.auto_bin_max=1024;
    option.per_instance=1;
    PC: coverpoint coverage_trans.PC;
    Imem_en: coverpoint coverage_trans.Imem_en;
    cmp_instr: coverpoint coverage_trans.cmp_instr;
    opcode: coverpoint coverage_trans.opcode;
    src1: coverpoint coverage_trans.src1;
    src2: coverpoint coverage_trans.src2;
    dest: coverpoint coverage_trans.dest;
    imm5: coverpoint coverage_trans.imm5;
    PCoffset9: coverpoint coverage_trans.PCoffset9;
    BaseR: coverpoint coverage_trans.BaseR;
    cnd_flags: coverpoint coverage_trans.cnd_flags;
    Instr_Dout: coverpoint coverage_trans.Instr_Dout;
    // pragma uvmf custom covergroup end
  endgroup

  covergroup alu_cg;

    // Cross for Register Adds 
    add_reg_cross : cross coverage_trans.src1,coverage_trans.src2,coverage_trans.dest,coverage_trans.opcode,coverage_trans.Instr_Dout[5]
      {
        bins all = add_reg_cross with (coverage_trans.Instr_Dout[5] == 0 && coverage_trans.opcode == 4'b0001 );
      }

    // Cross for Add immediates
    add_imm_cross : cross coverage_trans.src1,coverage_trans.imm5,coverage_trans.dest,coverage_trans.opcode,coverage_trans.Instr_Dout[5]
      {
        bins all = add_reg_cross with (coverage_trans.Instr_Dout[5] == 1 && coverage_trans.opcode == 4'b0001 );
      }
  endgroup

  // ****************************************************************************
  // FUNCTION : new()
  // This function is the standard SystemVerilog constructor.
  //
  function new(string name="", uvm_component parent=null);
    super.new(name,parent);
    instruction_memory_transaction_cg=new;
    `uvm_warning("COVERAGE_MODEL_REVIEW", "A covergroup has been constructed which may need review because of either generation or re-generation with merging.  Please note that transaction variables added as a result of re-generation and merging are not automatically added to the covergroup.  Remove this warning after the covergroup has been reviewed.")
  endfunction

  // ****************************************************************************
  // FUNCTION : build_phase()
  // This function is the standard UVM build_phase.
  //
  function void build_phase(uvm_phase phase);
    instruction_memory_transaction_cg.set_inst_name($sformatf("instruction_memory_transaction_cg_%s",get_full_name()));
  endfunction

  // ****************************************************************************
  // FUNCTION: write (T t)
  // This function is automatically executed when a transaction arrives on the
  // analysis_export.  It copies values from the variables in the transaction 
  // to local variables used to collect functional coverage.  
  //
  virtual function void write (T t);
    `uvm_info("COV","Received transaction",UVM_HIGH);
    coverage_trans = t;
    instruction_memory_transaction_cg.sample();
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

