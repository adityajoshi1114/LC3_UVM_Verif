//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This interface performs the instruction_memory signal monitoring.
//      It is accessed by the uvm instruction_memory monitor through a virtual
//      interface handle in the instruction_memory configuration.  It monitors the
//      signals passed in through the port connection named bus of
//      type instruction_memory_if.
//
//     Input signals from the instruction_memory_if are assigned to an internal input
//     signal with a _i suffix.  The _i signal should be used for sampling.
//
//     The input signal connections are as follows:
//       bus.signal -> signal_i 
//
//      Interface functions and tasks used by UVM components:
//             monitor(inout TRANS_T txn);
//                   This task receives the transaction, txn, from the
//                   UVM monitor and then populates variables in txn
//                   from values observed on bus activity.  This task
//                   blocks until an operation on the instruction_memory bus is complete.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
import uvmf_base_pkg_hdl::*;
import instruction_memory_pkg_hdl::*;
import instruction_memory_pkg::*;


interface instruction_memory_monitor_bfm 
  ( instruction_memory_if  bus );

`ifndef XRTL
// This code is to aid in debugging parameter mismatches between the BFM and its corresponding agent.
// Enable this debug by setting UVM_VERBOSITY to UVM_DEBUG
// Setting UVM_VERBOSITY to UVM_DEBUG causes all BFM's and all agents to display their parameter settings.
// All of the messages from this feature have a UVM messaging id value of "CFG"
// The transcript or run.log can be parsed to ensure BFM parameter settings match its corresponding agents parameter settings.
import uvm_pkg::*;
`include "uvm_macros.svh"
initial begin : bfm_vs_agent_parameter_debug
  `uvm_info("CFG", 
      $psprintf("The BFM at '%m' has the following parameters: ", ),
      UVM_DEBUG)
end
`endif


 instruction_memory_transaction  
                      monitored_trans;
 

  // Config value to determine if this is an initiator or a responder 
  uvmf_initiator_responder_t initiator_responder;
  // Custom configuration variables.  
  // These are set using the configure function which is called during the UVM connect_phase

  tri clock_i;
  tri reset_i;
  tri [15:0] PC_i;
  tri  instrmem_rd_i;
  tri [15:0] instr_dout_i;
  tri  complete_instr_i;
  assign clock_i = bus.clock;
  assign reset_i = bus.reset;
  assign PC_i = bus.PC;
  assign instrmem_rd_i = bus.instrmem_rd;
  assign instr_dout_i = bus.instr_dout;
  assign complete_instr_i = bus.complete_instr;

  // Proxy handle to UVM monitor
  instruction_memory_pkg::instruction_memory_monitor  proxy;

  // pragma uvmf custom interface_item_additional begin
  // pragma uvmf custom interface_item_additional end
  
  //******************************************************************                         
  task wait_for_reset(); 
    @(posedge clock_i) ;                                                                    
    do_wait_for_reset();                                                                   
  endtask                                                                                   

  // ****************************************************************************              
  task do_wait_for_reset(); 
  // pragma uvmf custom reset_condition begin
    wait ( reset_i === 0 ) ;                                                                   
  // pragma uvmf custom reset_condition end                                                                
  endtask    

  //******************************************************************                         
 
  task wait_for_num_clocks(input int unsigned count); 
    @(posedge clock_i);  
                                                                   
    repeat (count-1) @(posedge clock_i);                                                    
  endtask      

  //******************************************************************                         
  event go;                                                                                 
  function void start_monitoring();  
    -> go;
  endfunction                                                                               
  
  // ****************************************************************************              
  initial begin                                                                             
    @go;                                                                                   
    forever begin                                                                        
      monitored_trans = new("monitored_trans");
      do_monitor( ); 
    end                                                                                    
  end                                                                                       

  //******************************************************************
  // The configure() function is used to pass agent configuration
  // variables to the monitor BFM.  It is called by the monitor within
  // the agent at the beginning of the simulation.  It may be called 
  // during the simulation if agent configuration variables are updated
  // and the monitor BFM needs to be aware of the new configuration 
  // variables.
  //
    function void configure(instruction_memory_configuration 
                          
                         instruction_memory_configuration_arg
                         );  
    initiator_responder = instruction_memory_configuration_arg.initiator_responder;
  // pragma uvmf custom configure begin
  // pragma uvmf custom configure end
  endfunction   


  // ****************************************************************************  
  task do_monitor();
    //
    // Available struct members:
    //     //    monitored_trans.PC
    //     //    monitored_trans.Imem_en
    //     //    monitored_trans.cmp_instr
    //     //    monitored_trans.opcode
    //     //    monitored_trans.src1
    //     //    monitored_trans.src2
    //     //    monitored_trans.dest
    //     //    monitored_trans.imm5
    //     //    monitored_trans.PCoffset9
    //     //    monitored_trans.BaseR
    //     //    monitored_trans.cnd_flags
    //     //    monitored_trans.Instr_Dout
    //     //
    // Reference code;
    //    How to wait for signal value
    //      while (control_signal === 1'b1) @(posedge clock_i);
    //    
    //    How to assign a transaction variable, named xyz, from a signal.   
    //    All available input signals listed.
    //      monitored_trans.xyz = PC_i;  //    [15:0] 
    //      monitored_trans.xyz = instrmem_rd_i;  //     
    //      monitored_trans.xyz = instr_dout_i;  //    [15:0] 
    //      monitored_trans.xyz = complete_instr_i;  //     
    // pragma uvmf custom do_monitor begin
    // UVMF_CHANGE_ME : Implement protocol monitoring.  The commented reference code 
    // below are examples of how to capture signal values and assign them to 
    // structure members.  All available input signals are listed.  The 'while' 
    // code example shows how to wait for a synchronous flow control signal.  This
    // task should return when a complete transfer has been observed.  Once this task is
    // exited with captured values, it is then called again to wait for and observe 
    // the next transfer. One clock cycle is consumed between calls to do_monitor.
    // First Transaction 
    if (reset_i === 1'b1) begin 
      do_wait_for_reset();
      @(posedge clock_i);
    end
    
    if (complete_instr_i == 0) begin // If a valid instruction has been sent this cycle
      @(posedge complete_instr_i);
      @(posedge clock_i);
    end
    finish_monitoring();
    // pragma uvmf custom do_monitor end
  endtask         

  task finish_monitoring();
    // To fix casting issues
    reg_t src1_bus, src2_bus, src_bus, dest_bus, BaseR_bus;
    nzp_t cnd_flags_bus;
    opcode_t opcode_bus;
    monitored_trans.start_time = $time;
    @(negedge clock_i);   // Capture values at negedge
    monitored_trans.PC  = PC_i;
    monitored_trans.Imem_en = instrmem_rd_i;
    monitored_trans.Instr_Dout  = instr_dout_i;
    if (!$cast(opcode_bus,instr_dout_i[15:12])) $fatal;
    if (!$cast(src1_bus,instr_dout_i[8:6])) $fatal;
    if (!$cast(src2_bus,instr_dout_i[2:0])) $fatal;
    if (!$cast(src_bus, instr_dout_i[11:9])) $fatal;
    if (!$cast(dest_bus,instr_dout_i[11:9])) $fatal;
    if (!$cast(BaseR_bus,instr_dout_i[8:6])) $fatal;
    if (instr_dout_i[11:9] != 3'b000) begin 
      if (!$cast(cnd_flags_bus,instr_dout_i[11:9])) $fatal;
    end
    monitored_trans.opcode = opcode_bus;
    monitored_trans.src1 = src1_bus ;
    monitored_trans.src2 = src2_bus ;
    monitored_trans.src  = src_bus ;
    monitored_trans.dest = dest_bus ;
    monitored_trans.imm5 = instr_dout_i[4:0];
    monitored_trans.PCoffset9 = instr_dout_i[8:0];
    monitored_trans.PCoffset6 = instr_dout_i[5:0];
    monitored_trans.BaseR = BaseR_bus;
    if (instr_dout_i[11:9] != 3'b000) begin 
      monitored_trans.cnd_flags = cnd_flags_bus;
    end
    monitored_trans.cmp_instr = complete_instr_i;
    @(posedge clock_i);   // Move to end of transaction
    monitored_trans.end_time = $time;
    proxy.notify_transaction( monitored_trans ); 
  endtask
  
 
endinterface

// pragma uvmf custom external begin
// pragma uvmf custom external end

